module hex(input [15:0] in,
           output reg [27:0] out);
    
    always @(*) begin
<<<<<<< Updated upstream
        case (in)
            16'h001D: out = ~28'h000035e;
            16'hF01d: out =  ~28'h00000f1;
            16'h0000: out =  ~28'h0000000;
            default: out =  ~28'hfffffff;
        endcase
=======
        case (in[3:0])
            4'b0000: out[6:0] = ~7'h3F;
            4'b0001: out[6:0] = ~7'h06;
            4'b0010: out[6:0] = ~7'h5B;
            4'b0011: out[6:0] = ~7'h4F;
            4'b0100: out[6:0] = ~7'h66;
            4'b0101: out[6:0] = ~7'h6D;
            4'b0110: out[6:0] = ~7'h7D;
            4'b0111: out[6:0] = ~7'h07;
            4'b1000: out[6:0] = ~7'h7F;
            4'b1001: out[6:0] = ~7'h6F;
            4'b1010: out[6:0] = ~7'h77;
            4'b1011: out[6:0] = ~7'h7C;
            4'b1100: out[6:0] = ~7'h39;
            4'b1101: out[6:0] = ~7'h5E;
            4'b1110: out[6:0] = ~7'h79;
            4'b1111: out[6:0] = ~7'h71;
        endcase
        case (in[7:4])
            4'b0000: out[13:7] = ~7'h3F;
            4'b0001: out[13:7] = ~7'h06;
            4'b0010: out[13:7] = ~7'h5B;
            4'b0011: out[13:7] = ~7'h4F;
            4'b0100: out[13:7] = ~7'h66;
            4'b0101: out[13:7] = ~7'h6D;
            4'b0110: out[13:7] = ~7'h7D;
            4'b0111: out[13:7] = ~7'h07;
            4'b1000: out[13:7] = ~7'h7F;
            4'b1001: out[13:7] = ~7'h6F;
            4'b1010: out[13:7] = ~7'h77;
            4'b1011: out[13:7] = ~7'h7C;
            4'b1100: out[13:7] = ~7'h39;
            4'b1101: out[13:7] = ~7'h5E;
            4'b1110: out[13:7] = ~7'h79;
            4'b1111: out[13:7] = ~7'h71;
        endcase
         case (in[11:8])
            4'b0000: out[20:14] = ~7'h3F;
            4'b0001: out[20:14] = ~7'h06;
            4'b0010: out[20:14] = ~7'h5B;
            4'b0011: out[20:14] = ~7'h4F;
            4'b0100: out[20:14] = ~7'h66;
            4'b0101: out[20:14] = ~7'h6D;
            4'b0110: out[20:14] = ~7'h7D;
            4'b0111: out[20:14] = ~7'h07;
            4'b1000: out[20:14] = ~7'h7F;
            4'b1001: out[20:14] = ~7'h6F;
            4'b1010: out[20:14] = ~7'h77;
            4'b1011: out[20:14] = ~7'h7C;
            4'b1100: out[20:14] = ~7'h39;
            4'b1101: out[20:14] = ~7'h5E;
            4'b1110: out[20:14] = ~7'h79;
            4'b1111: out[20:14] = ~7'h71;
        endcase
         case (in[15:12])
            4'b0000: out[27:21] = ~7'h3F;
            4'b0001: out[27:21] = ~7'h06;
            4'b0010: out[27:21] = ~7'h5B;
            4'b0011: out[27:21] = ~7'h4F;
            4'b0100: out[27:21] = ~7'h66;
            4'b0101: out[27:21] = ~7'h6D;
            4'b0110: out[27:21] = ~7'h7D;
            4'b0111: out[27:21] = ~7'h07;
            4'b1000: out[27:21] = ~7'h7F;
            4'b1001: out[27:21] = ~7'h6F;
            4'b1010: out[27:21] = ~7'h77;
            4'b1011: out[27:21] = ~7'h7C;
            4'b1100: out[27:21] = ~7'h39;
            4'b1101: out[27:21] = ~7'h5E;
            4'b1110: out[27:21] = ~7'h79;
            4'b1111: out[27:21] = ~7'h71;
        endcase
>>>>>>> Stashed changes
    end
    
endmodule
